import PAClib :: *;

import Controller :: *;
import DataTypes :: *;
import Headers :: *;
import SpecialFIFOF :: *;
import Settings :: *;
import RetryHandleSQ :: *;
import ReqGenSQ :: *;
import RespHandleSQ :: *;
import WorkCompGenSQ :: *;
import Utils :: *;

interface SQ;
    interface DataStreamPipeOut rdmaReqDataStreamPipeOut;
    interface PipeOut#(WorkComp) workCompPipeOut;
endinterface

module mkSQ#(
    Controller cntrl,
    PipeOut#(WorkReq) workReqPipeIn,
    DmaReadSrv dmaReadSrv,
    DmaWriteSrv dmaWriteSrv,
    DataStreamPipeOut rdmaRespPipeIn,
    PipeOut#(WorkCompStatus) workCompStatusPipeInFromRQ
)(SQ);
    PendingWorkReqBuf pendingWorkReqBuf <- mkScanFIFOF;

    let newPendingWorkReqPipeOut <- mkNewPendingWorkReqPipeOut(workReqPipeIn);
    // let retryPendingWorkReqPipeOut = scanQ2PipeOut(pendingWorkReqScan);

    let retryHandler <- mkRetryHandleSQ(cntrl, pendingWorkReqBuf.scanIfc);
    let notRetrying = retryHandler.isRetryDone;

    let pendingWorkReqPipeOut = muxPipeOut(
        notRetrying,
        newPendingWorkReqPipeOut,
        retryHandler.retryWorkReqPipeOut
    );
    let reqGenSQ <- mkReqGenSQ(
        cntrl, dmaReadSrv, pendingWorkReqPipeOut, pendingWorkReqBuf.fifoIfc.notEmpty
    );

    let headerAndMetaDataAndPayloadPipeOut <- mkExtractHeaderFromRdmaPktPipeOut(
        rdmaRespPipeIn
    );
    let pktMetaDataAndPayloadPipeOut <- mkInputRdmaPktBufAndHeaderValidation(
        headerAndMetaDataAndPayloadPipeOut, cntrl.getPMTU
    );

    let respHandleSQ <- mkRespHandleSQ(
        cntrl,
        convertFifo2PipeOut(pendingWorkReqBuf.fifoIfc),
        pktMetaDataAndPayloadPipeOut.pktMetaData,
        retryHandler
    );

    let payloadConsumer <- mkPayloadConsumer(
        cntrl,
        pktMetaDataAndPayloadPipeOut.payload,
        dmaWriteSrv,
        respHandleSQ.payloadConReqPipeOut
    );

    let wcPipeOut <- mkWorkCompGenSQ(
        cntrl,
        payloadConsumer.respPipeOut,
        reqGenSQ.workCompGenReqPipeOut,
        respHandleSQ.workCompGenReqPipeOut,
        workCompStatusPipeInFromRQ
    );

    interface rdmaReqDataStreamPipeOut = reqGenSQ.rdmaReqDataStreamPipeOut;
    interface workCompPipeOut = wcPipeOut;
endmodule

interface RQ;
    interface DataStreamPipeOut rdmaRespDataStreamPipeOut;
    interface WorkCompGenRQ wcGenRQ;
endinterface

module mkRQ#(
    Controller cntrl,
    DmaReadSrv dmaReadSrv,
    DmaWriteSrv dmaWriteSrv,
    DataStreamPipeOut payloadPipeIn,
    PermCheckMR permCheckMR,
    RecvReqBuf recvReqBuf,
    PipeOut#(RdmaPktMetaData) pktMetaDataPipeIn
)(ReqHandleRQ);
    let payloadGenerator <- mkPayloadGenerator(
        cntrl, dmaReadSrv, convertFifo2PipeOut(payloadGenReqOutQ)
    );
    let dupReadAtomicCache <- mkDupReadAtomicCache(cntrl);

    let reqHandlerRQ <- mkReqHandleRQ(
        cntrl,
        dmaReadSrv,
        permCheckMR,
        dupReadAtomicCache,
        recvReqBuf,
        pktMetaDataPipeIn
    );

    let payloadConsumer <- mkPayloadConsumer(
        cntrl,
        payloadPipeIn,
        dmaWriteSrv,
        reqHandlerRQ.payloadConReqPipeOut
    );

    let workCompGenRQ <- mkWorkCompGenRQ(
        cntrl,
        payloadConsumer.respPipeOut,
        reqHandlerRQ.workCompGenReqPipeOut
    );

    interface rdmaRespDataStreamPipeOut = reqHandlerRQ.rdmaRespDataStreamPipeOut;
    interface wcGenRQ = workCompGenRQ;
endmodule

interface QP;
    PipeOut#(WorkComp) workCompPipeOutSQ;
    PipeOut#(WorkComp) workCompPipeOutRQ;
endinterface

module mkQP#()(QP);
    // TODO: if WR queue is empty, then error flush is done
    if (!workReqPipeIn.notEmpty) begin
        // Notify controller when flush done
        cntrl.errFlushDone;
        $display(
            "time=%0d: error flush done, pendingWorkCompQ4SQ.notEmpty=",
            $time, fshow(pendingWorkCompQ4SQ.notEmpty)
        );
    end
endmodule
